// Copyright 2025 Maktab-e-Digital Systems Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description:
//    Header file containing localparam definitions for Y (Luma) Huffman encoding.
//    These parameters define the DC and AC Huffman code lengths and codes,
//    as well as the AC run-length Huffman mapping.
//
// Author:Rameen
// Date:15th July,2025.

`ifndef CB_HUFF_CONSTANTS_SVH
`define CB_HUFF_CONSTANTS_SVH

localparam int Cb_DC_code_length [0:11] = '{
    2, 2, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11
};

localparam logic [10:0] Cb_DC [0:11] = '{
    11'b00000000000,
    11'b01000000000,
    11'b10000000000,
    11'b11000000000,
    11'b11100000000,
    11'b11110000000,
    11'b11111000000,
    11'b11111100000,
    11'b11111110000,
    11'b11111111000,
    11'b11111111100,
    11'b11111111110
};

localparam int Cb_AC_code_length [0:161] = '{
    // 0 - 35: Explicit values
    2, 2, 3, 4, 4, 4, 5, 5, 5, 6, 6, 7, 7, 7, 7,
    8, 8, 8, 9, 9, 9, 9, 9, 10, 10, 10, 10, 10,
    11, 11, 11, 11, 12, 12, 12, 12,
    
    // 36 - 161: Repeated value = 16
    {126{16}}
};

localparam logic [15:0] Cb_AC [0:161] = '{
  16'h0000, 16'h4000, 16'h8000, 16'hA000, 16'hB000, 16'hC000, 16'hD000, 16'hD800,
  16'hE000, 16'hE800, 16'hEC00, 16'hF000, 16'hF200, 16'hF400, 16'hF600, 16'hF800,
  16'hF900, 16'hFA00, 16'hFB00, 16'hFB80, 16'hFC00, 16'hFC80, 16'hFD00, 16'hFD80,
  16'hFDC0, 16'hFE00, 16'hFE40, 16'hFE80, 16'hFEC0, 16'hFEE0, 16'hFF00, 16'hFF20,
  16'hFF40, 16'hFF50, 16'hFF60, 16'hFF70, 16'hFF80, 16'hFF82, 16'hFF83, 16'hFF84,
  16'hFF85, 16'hFF86, 16'hFF87, 16'hFF88, 16'hFF89, 16'hFF8A, 16'hFF8B, 16'hFF8C,
  16'hFF8D, 16'hFF8E, 16'hFF8F, 16'hFF90, 16'hFF91, 16'hFF92, 16'hFF93, 16'hFF94,
  16'hFF95, 16'hFF96, 16'hFF97, 16'hFF98, 16'hFF99, 16'hFF9A, 16'hFF9B, 16'hFF9C,
  16'hFF9D, 16'hFF9E, 16'hFF9F, 16'hFFA0, 16'hFFA1, 16'hFFA2, 16'hFFA3, 16'hFFA4,
  16'hFFA5, 16'hFFA6, 16'hFFA7, 16'hFFA8, 16'hFFA9, 16'hFFAA, 16'hFFAB, 16'hFFAC,
  16'hFFAD, 16'hFFAE, 16'hFFAF, 16'hFFB0, 16'hFFB1, 16'hFFB2, 16'hFFB3, 16'hFFB4,
  16'hFFB5, 16'hFFB6, 16'hFFB7, 16'hFFB8, 16'hFFB9, 16'hFFBA, 16'hFFBB, 16'hFFBC,
  16'hFFBD, 16'hFFBE, 16'hFFBF, 16'hFFC0, 16'hFFC1, 16'hFFC2, 16'hFFC3, 16'hFFC4,
  16'hFFC5, 16'hFFC6, 16'hFFC7, 16'hFFC8, 16'hFFC9, 16'hFFCA, 16'hFFCB, 16'hFFCC,
  16'hFFCD, 16'hFFCE, 16'hFFCF, 16'hFFD0, 16'hFFD1, 16'hFFD2, 16'hFFD3, 16'hFFD4,
  16'hFFD5, 16'hFFD6, 16'hFFD7, 16'hFFD8, 16'hFFD9, 16'hFFDA, 16'hFFDB, 16'hFFDC,
  16'hFFDD, 16'hFFDE, 16'hFFDF, 16'hFFE0, 16'hFFE1, 16'hFFE2, 16'hFFE3, 16'hFFE4,
  16'hFFE5, 16'hFFE6, 16'hFFE7, 16'hFFE8, 16'hFFE9, 16'hFFEA, 16'hFFEB, 16'hFFEC,
  16'hFFED, 16'hFFEE, 16'hFFEF, 16'hFFF0, 16'hFFF1, 16'hFFF2, 16'hFFF3, 16'hFFF4,
  16'hFFF5, 16'hFFF6, 16'hFFF7, 16'hFFF8, 16'hFFF9, 16'hFFFA, 16'hFFFB, 16'hFFFC,
  16'hFFFD, 16'hFFFE
};

localparam int Cb_AC_run_code [0:250] = '{
  3, // [0]
  0, // [1]
  1, // [2]
  2, // [3]
  4, // [4]
  6, // [5]
  11, // [6]
  15, // [7]
  23, // [8]
  37, // [9]
  38, // [10]
  0, // [11–15] default
  0, // [16]
  5, // [17]
  7, // [18]
  12, // [19]
  18, // [20]
  28, // [21]
  39, // [22]
  40, // [23]
  41, // [24]
  42, // [25]
  43, // [26]
  0, // [27–31]
  0, // [32]
  8, // [33]
  16, // [34]
  24, // [35]
  32, // [36]
  44, // [37]
  45, // [38]
  46, // [39]
  47, // [40]
  48, // [41]
  49, // [42]
  0,  // [43]
  50, // [52]
  51, // [53]
  52, // [54]
  53, // [55]
  54, // [56]
  55, // [57]
  56, // [58]
  0, // [59–63]
  0, // [64]
  25, // [65]
  57, // [66]
  59, // [67]
  58, // [68]
  59, // [69]
  60, // [70]
  61, // [71]
  62, // [72]
  63, // [73]
  64, // [74]
  0,  // [75–79]
  13, // [81]
  29, // [82]
  65, // [83]
  66, // [84]
  67, // [85]
  68, // [86]
  69, // [87]
  70, // [88]
  71, // [89]
  72, // [90]
  0,  // [91–95]
  14, // [97]
  34, // [98]
  73, // [99]
  74, // [100]
  75, // [101]
  76, // [102]
  77, // [103]
  78, // [104]
  79, // [105]
  80, // [106]
  0,  // [107–111]
  17, // [113]
  81, // [114]
  81, // [115]
  82, // [116]
  83, // [117]
  84, // [118]
  85, // [119]
  86, // [120]
  87, // [121]
  88, // [122]
  0,  // [123–127]
  10, // [128]
  89, // [131]
  90, // [132]
  91, // [133]
  92, // [134]
  93, // [135]
  94, // [136]
  95, // [137]
  96, // [138]
  0,  // [139–143]
  21, // [145]
  97, // [146]
  98, // [147]
  99, // [148]
 100, // [149]
 101, // [150]
 102, // [151]
 103, // [152]
 104, // [153]
 105, // [154]
  0,  // [155–161]
 106, // [162]
 107, // [163]
 108, // [164]
 109, // [165]
 110, // [166]
 111, // [167]
 112, // [168]
 113, // [169]
 114, // [170]
  0,  // [171–176]
  26, // [177]
 115, // [178]
 116, // [179]
 117, // [180]
 118, // [181]
 119, // [182]
 120, // [183]
 121, // [184]
 122, // [185]
 123, // [186]
  0,  // [187–192]
  27, // [193]
 124, // [194]
 125, // [195]
 126, // [196]
 127, // [197]
 128, // [198]
 129, // [199]
 130, // [200]
 131, // [201]
 132, // [202]
  0,  // [203–208]
  30, // [209]
 133, // [210]
 134, // [211]
 135, // [212]
 136, // [213]
 137, // [214]
 138, // [215]
 139, // [216]
 140, // [217]
 141, // [218]
  0,  // [219–224]
 142, // [225]
 143, // [226]
 144, // [227]
 145, // [228]
 146, // [229]
 147, // [230]
 148, // [231]
 149, // [232]
 150, // [233]
 151, // [234]
  0,  // [235–240]
 152, // [241]
 153, // [242]
 154, // [243]
 155, // [244]
 156, // [245]
 157, // [246]
 158, // [247]
 159, // [248]
 160, // [249]
 161  // [250]
};
`endif
